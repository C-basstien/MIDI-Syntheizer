library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;




entity MIDI_ROM is
  port
  (
  	rom_fsm_address  : 	in  std_logic_vector(9 downto 0);
  	rom_comp_address :	in  std_logic_vector(9 downto 0);
  	rom_vlq_address  : 	in  std_logic_vector(9 downto 0);
  
  	rom_fsm_out    : 	out std_logic_vector(7 downto 0);
  	rom_comp_out    : 	out std_logic_vector(7 downto 0);
  	rom_vlq_out    : 	out std_logic_vector(7 downto 0);
  	
  );
end ROM;

architecture MIDI_ROM_A of MIDI_ROM is
  type     tab_rom is array (0 to 567) of std_logic_vector(7 downto 0);
  constant filter_rom : tab_rom := -- Tableau des coefficients du filtre
    (
		0 => "01001101" , 1 => "01010100" , 2 => "01101000" , 3 => "01100100" , 
		4 => "00000000" , 5 => "00000000" , 6 => "00000000" , 7 => "00000110" , 
		8 => "00000000" , 9 => "00000001" , 10 => "00000000" , 11 => "00000010" , 
		12 => "00000011" , 13 => "11000000" , 14 => "01001101" , 15 => "01010100" , 
		16 => "01110010" , 17 => "01101011" , 18 => "00000000" , 19 => "00000000" , 
		20 => "00000000" , 21 => "00011001" , 22 => "00000000" , 23 => "11111111" , 
		24 => "01011000" , 25 => "00000100" , 26 => "00000100" , 27 => "00000010" , 
		28 => "00011000" , 29 => "00001000" , 30 => "00000000" , 31 => "11111111" , 
		32 => "01011001" , 33 => "00000010" , 34 => "00000000" , 35 => "00000000" , 
		36 => "00000000" , 37 => "11111111" , 38 => "01010001" , 39 => "00000011" , 
		40 => "00001001" , 41 => "00100111" , 42 => "11000000" , 43 => "00000001" , 
		44 => "11111111" , 45 => "00101111" , 46 => "00000000" , 47 => "01001101" , 
		48 => "01010100" , 49 => "01110010" , 50 => "01101011" , 51 => "00000000" , 
		52 => "00000000" , 53 => "00000001" , 54 => "11111111" , 55 => "00000000" , 
		56 => "11000000" , 57 => "00000000" , 58 => "00000000" , 59 => "10110000" , 
		60 => "01111001" , 61 => "00000000" , 62 => "00000000" , 63 => "10110000" , 
		64 => "01000000" , 65 => "00000000" , 66 => "00000000" , 67 => "10110000" , 
		68 => "01011011" , 69 => "00110000" , 70 => "00000000" , 71 => "10110000" , 
		72 => "00001010" , 73 => "00110011" , 74 => "00000000" , 75 => "10110000" , 
		76 => "00000111" , 77 => "01100100" , 78 => "00000000" , 79 => "10010000" , 
		80 => "00111100" , 81 => "01000101" , 82 => "00000000" , 83 => "10110000" , 
		84 => "01111001" , 85 => "00000000" , 86 => "00000000" , 87 => "10110000" , 
		88 => "01000000" , 89 => "00000000" , 90 => "00000000" , 91 => "10110000" , 
		92 => "01011011" , 93 => "00110000" , 94 => "00000000" , 95 => "10110000" , 
		96 => "00001010" , 97 => "00110011" , 98 => "00000000" , 99 => "10110000" , 
		100 => "00000111" , 101 => "01100100" , 102 => "00000000" , 103 => "11111111" , 
		104 => "00000011" , 105 => "00000101" , 106 => "01010000" , 107 => "01101001" , 
		108 => "01100001" , 109 => "01101110" , 110 => "01101111" , 111 => "00000000" , 
		112 => "10010000" , 113 => "00110000" , 114 => "01001010" , 115 => "10000111" , 
		116 => "01000000" , 117 => "10000000" , 118 => "00111100" , 119 => "00000000" , 
		120 => "00000000" , 121 => "10010000" , 122 => "00111100" , 123 => "01001100" , 
		124 => "00000000" , 125 => "10000000" , 126 => "00110000" , 127 => "00000000" , 
		128 => "00000000" , 129 => "10010000" , 130 => "00110111" , 131 => "01001111" , 
		132 => "10000111" , 133 => "01000000" , 134 => "10000000" , 135 => "00111100" , 
		136 => "00000000" , 137 => "00000000" , 138 => "10010000" , 139 => "00111100" , 
		140 => "01001010" , 141 => "00000000" , 142 => "10000000" , 143 => "00110111" , 
		144 => "00000000" , 145 => "00000000" , 146 => "10010000" , 147 => "00110100" , 
		148 => "01001001" , 149 => "10000111" , 150 => "01000000" , 151 => "10000000" , 
		152 => "00111100" , 153 => "00000000" , 154 => "00000000" , 155 => "10010000" , 
		156 => "00111110" , 157 => "01010000" , 158 => "00000000" , 159 => "10000000" , 
		160 => "00110100" , 161 => "00000000" , 162 => "00000000" , 163 => "10010000" , 
		164 => "00110111" , 165 => "01001101" , 166 => "10000111" , 167 => "01000000" , 
		168 => "10000000" , 169 => "00111110" , 170 => "00000000" , 171 => "00000000" , 
		172 => "10010000" , 173 => "01000000" , 174 => "01010000" , 175 => "00000000" , 
		176 => "10000000" , 177 => "00110111" , 178 => "00000000" , 179 => "00000000" , 
		180 => "10010000" , 181 => "00110000" , 182 => "01001001" , 183 => "10000111" , 
		184 => "01000000" , 185 => "10000000" , 186 => "00110000" , 187 => "00000000" , 
		188 => "00000000" , 189 => "10010000" , 190 => "00110111" , 191 => "01010001" , 
		192 => "10000111" , 193 => "01000000" , 194 => "10000000" , 195 => "01000000" , 
		196 => "00000000" , 197 => "00000000" , 198 => "10010000" , 199 => "00111110" , 
		200 => "01000111" , 201 => "00000000" , 202 => "10000000" , 203 => "00110111" , 
		204 => "00000000" , 205 => "00000000" , 206 => "10010000" , 207 => "00110101" , 
		208 => "01001001" , 209 => "10000111" , 210 => "01000000" , 211 => "10000000" , 
		212 => "00110101" , 213 => "00000000" , 214 => "00000000" , 215 => "10010000" , 
		216 => "00110111" , 217 => "01001110" , 218 => "10000111" , 219 => "01000000" , 
		220 => "10000000" , 221 => "00111110" , 222 => "00000000" , 223 => "00000000" , 
		224 => "10010000" , 225 => "00111100" , 226 => "01000111" , 227 => "00000000" , 
		228 => "10000000" , 229 => "00110111" , 230 => "00000000" , 231 => "00000000" , 
		232 => "10010000" , 233 => "00110100" , 234 => "01010001" , 235 => "10000111" , 
		236 => "01000000" , 237 => "10000000" , 238 => "00111100" , 239 => "00000000" , 
		240 => "00000000" , 241 => "10010000" , 242 => "01000000" , 243 => "01010010" , 
		244 => "00000000" , 245 => "10000000" , 246 => "00110100" , 247 => "00000000" , 
		248 => "00000000" , 249 => "10010000" , 250 => "00110111" , 251 => "01010010" , 
		252 => "10000111" , 253 => "01000000" , 254 => "10000000" , 255 => "01000000" , 
		256 => "00000000" , 257 => "00000000" , 258 => "10010000" , 259 => "00111110" , 
		260 => "01001110" , 261 => "00000000" , 262 => "10000000" , 263 => "00110111" , 
		264 => "00000000" , 265 => "00000000" , 266 => "10010000" , 267 => "00110101" , 
		268 => "01000111" , 269 => "10000111" , 270 => "01000000" , 271 => "10000000" , 
		272 => "00111110" , 273 => "00000000" , 274 => "00000000" , 275 => "10010000" , 
		276 => "00111110" , 277 => "01010001" , 278 => "00000000" , 279 => "10000000" , 
		280 => "00110101" , 281 => "00000000" , 282 => "00000000" , 283 => "10010000" , 
		284 => "00110010" , 285 => "01000110" , 286 => "10000111" , 287 => "01000000" , 
		288 => "10000000" , 289 => "00111110" , 290 => "00000000" , 291 => "00000000" , 
		292 => "10010000" , 293 => "00111100" , 294 => "01000101" , 295 => "00000000" , 
		296 => "10000000" , 297 => "00110010" , 298 => "00000000" , 299 => "00000000" , 
		300 => "10010000" , 301 => "00110100" , 302 => "01001110" , 303 => "10000111" , 
		304 => "01000000" , 305 => "10000000" , 306 => "00110100" , 307 => "00000000" , 
		308 => "00000000" , 309 => "10010000" , 310 => "00110111" , 311 => "01001101" , 
		312 => "10000111" , 313 => "01000000" , 314 => "10000000" , 315 => "00110111" , 
		316 => "00000000" , 317 => "00000000" , 318 => "10010000" , 319 => "00110101" , 
		320 => "01001010" , 321 => "10000111" , 322 => "01000000" , 323 => "10000000" , 
		324 => "00110101" , 325 => "00000000" , 326 => "00000000" , 327 => "10010000" , 
		328 => "00110010" , 329 => "01000111" , 330 => "10000111" , 331 => "01000000" , 
		332 => "10000000" , 333 => "00111100" , 334 => "00000000" , 335 => "00000000" , 
		336 => "10010000" , 337 => "00111100" , 338 => "01001101" , 339 => "00000000" , 
		340 => "10000000" , 341 => "00110010" , 342 => "00000000" , 343 => "00000000" , 
		344 => "10010000" , 345 => "00110000" , 346 => "01001000" , 347 => "10000111" , 
		348 => "01000000" , 349 => "10000000" , 350 => "00111100" , 351 => "00000000" , 
		352 => "00000000" , 353 => "10010000" , 354 => "00111100" , 355 => "01001010" , 
		356 => "00000000" , 357 => "10000000" , 358 => "00110000" , 359 => "00000000" , 
		360 => "00000000" , 361 => "10010000" , 362 => "00110111" , 363 => "01010010" , 
		364 => "10000111" , 365 => "01000000" , 366 => "10000000" , 367 => "00111100" , 
		368 => "00000000" , 369 => "00000000" , 370 => "10010000" , 371 => "00111100" , 
		372 => "01001101" , 373 => "00000000" , 374 => "10000000" , 375 => "00110111" , 
		376 => "00000000" , 377 => "00000000" , 378 => "10010000" , 379 => "00110100" , 
		380 => "01001100" , 381 => "10000111" , 382 => "01000000" , 383 => "10000000" , 
		384 => "00111100" , 385 => "00000000" , 386 => "00000000" , 387 => "10010000" , 
		388 => "00111110" , 389 => "01010001" , 390 => "00000000" , 391 => "10000000" , 
		392 => "00110100" , 393 => "00000000" , 394 => "00000000" , 395 => "10010000" , 
		396 => "00110111" , 397 => "01010001" , 398 => "10000111" , 399 => "01000000" , 
		400 => "10000000" , 401 => "00111110" , 402 => "00000000" , 403 => "00000000" , 
		404 => "10010000" , 405 => "01000000" , 406 => "01010011" , 407 => "00000000" , 
		408 => "10000000" , 409 => "00110111" , 410 => "00000000" , 411 => "00000000" , 
		412 => "10010000" , 413 => "00110000" , 414 => "01000110" , 415 => "10000111" , 
		416 => "01000000" , 417 => "10000000" , 418 => "00110000" , 419 => "00000000" , 
		420 => "00000000" , 421 => "10010000" , 422 => "00110111" , 423 => "01010010" , 
		424 => "10000111" , 425 => "01000000" , 426 => "10000000" , 427 => "01000000" , 
		428 => "00000000" , 429 => "00000000" , 430 => "10010000" , 431 => "00111110" , 
		432 => "01001000" , 433 => "00000000" , 434 => "10000000" , 435 => "00110111" , 
		436 => "00000000" , 437 => "00000000" , 438 => "10010000" , 439 => "00110101" , 
		440 => "01001010" , 441 => "10000111" , 442 => "01000000" , 443 => "10000000" , 
		444 => "00110101" , 445 => "00000000" , 446 => "00000000" , 447 => "10010000" , 
		448 => "00110111" , 449 => "01001111" , 450 => "10000111" , 451 => "01000000" , 
		452 => "10000000" , 453 => "00111110" , 454 => "00000000" , 455 => "00000000" , 
		456 => "10010000" , 457 => "00111100" , 458 => "01001000" , 459 => "00000000" , 
		460 => "10000000" , 461 => "00110111" , 462 => "00000000" , 463 => "00000000" , 
		464 => "10010000" , 465 => "00110100" , 466 => "01000111" , 467 => "10000111" , 
		468 => "01000000" , 469 => "10000000" , 470 => "00111100" , 471 => "00000000" , 
		472 => "00000000" , 473 => "10010000" , 474 => "01000000" , 475 => "01010111" , 
		476 => "00000000" , 477 => "10000000" , 478 => "00110100" , 479 => "00000000" , 
		480 => "00000000" , 481 => "10010000" , 482 => "00110111" , 483 => "01001110" , 
		484 => "10000111" , 485 => "01000000" , 486 => "10000000" , 487 => "01000000" , 
		488 => "00000000" , 489 => "00000000" , 490 => "10010000" , 491 => "00111110" , 
		492 => "01000100" , 493 => "00000000" , 494 => "10000000" , 495 => "00110111" , 
		496 => "00000000" , 497 => "00000000" , 498 => "10010000" , 499 => "00110101" , 
		500 => "01000111" , 501 => "10000111" , 502 => "01000000" , 503 => "10000000" , 
		504 => "00111110" , 505 => "00000000" , 506 => "00000000" , 507 => "10010000" , 
		508 => "00111110" , 509 => "01001011" , 510 => "00000000" , 511 => "10000000" , 
		512 => "00110101" , 513 => "00000000" , 514 => "00000000" , 515 => "10010000" , 
		516 => "00101111" , 517 => "01000110" , 518 => "10000111" , 519 => "01000000" , 
		520 => "10000000" , 521 => "00111110" , 522 => "00000000" , 523 => "00000000" , 
		524 => "10010000" , 525 => "00111100" , 526 => "01001000" , 527 => "00000000" , 
		528 => "10000000" , 529 => "00101111" , 530 => "00000000" , 531 => "00000000" , 
		532 => "10010000" , 533 => "00110000" , 534 => "01010010" , 535 => "10000111" , 
		536 => "01000000" , 537 => "10000000" , 538 => "00110000" , 539 => "00000000" , 
		540 => "00000000" , 541 => "10010000" , 542 => "00110111" , 543 => "01010101" , 
		544 => "10000111" , 545 => "01000000" , 546 => "10000000" , 547 => "00110111" , 
		548 => "00000000" , 549 => "00000000" , 550 => "10010000" , 551 => "00110000" , 
		552 => "01000110" , 553 => "10001111" , 554 => "00000000" , 555 => "10000000" , 
		556 => "00111100" , 557 => "00000000" , 558 => "00000000" , 559 => "10000000" , 
		560 => "00110000" , 561 => "00000000" , 562 => "00000001" , 563 => "11111111" , 
		564 => "00101111" , 565 => "00000000" , 566 => "11111111" , 567 => "11111111" 
	) ;

begin

  rom__fsm_out  <= filter_rom(to_integer(unsigned(rom_fsm_address))); --  valeur du coefficient demandé par la fsm
  rom_comp_out <= filter_rom(to_integer(unsigned(rom_comp_address))); -- valeur du coefficient demandé par le comparateur;
  rom_vlq_out  <= filter_rom(to_integer(unsigned(rom_vlq_address))); -- valeur du coefficient demandé par le calculateur de vlq
  

end A;
